En svart katt .
En gul fågel .
En vit elefant .
